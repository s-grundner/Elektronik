-- VHDL

/* [1.5 - 1] Which of the following are valid VHDL basic identifiers? Which are reserved words? 
 * Of the invalid identifiers, why are they invalid?
 * last_item 	-> valid
 * prev item 	-> invalid, contains space
 * value-1 		-> invalid, '-' is a special symbol
 * buffer 		-> invalid, is vhdl keyword
 * element#5 	-> invalid, '#' is a special symbol
 * _control		-> invalid, does not start with alphabetical character
 * 93_999		-> invalid, does not start with alphabetical character
 * entry_		-> valid
 */
 
/* [1.5 - 2] Rewrite the following decimal literals as hexadecimal literals.
 * 1		16#1#
 * 34		16#22#
 * 256.0	16#FF#
 * 0.5		16#0.8#
 */
 
/* [1.5 - 3] What decimal numbers are represented by the following literals?
 * 8#14#			12
 * 2#1000_0100# 	132
 * 6#2C#			44
 * 2.5E5			250_000
 * 2#1#E15			32_768
 * 2#0.101#			0.625
 */
 
/* [1.5 - 4] What is the difference between the literals
 * 16#23DF# = B#10_0011_1101_1111#
 * X"23DF" = B"0010_0011_1101_1111"
 */
 
 